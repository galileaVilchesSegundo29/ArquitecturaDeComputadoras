LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY or00 IS
    PORT(
        Ao, Bo: IN STD_LOGIC;
        Yo: OUT STD_LOGIC);
END or00;

ARCHITECTURE A_or00 OF or00 IS
BEGIN
    Yo <= Ao OR Bo;
END A_or00;