LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
USE PACKAGEALU00.ALL;

ENTITY TOPALU00 IS
PORT(
		CLK00: INOUT STD_LOGIC;
		ENABLE0:IN STD_LOGIC;
		CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		FUNCT0: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		INREGRS0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		INREGRT0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTALU0: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTFLAGINST0: INOUT STD_LOGIC;
		OUTFLAGAC0: INOUT STD_LOGIC		
	);
END TOPALU00;

ARCHITECTURE A_TOPALU00 OF TOPALU00 IS
SIGNAL SDATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN

	AL00: TOPDIV00 PORT MAP(CLK0 => CLK00,
							CDIV0 => CDIV00
							);
	
	AL01: ANDA00 PORT MAP(CLKA => CLK00,
							INFLAGA => OUTFLAGAC0,
							FUNCTA => FUNCT0,
							INRSA =>  INREGRS0,
							INRTA  => INREGRT0,
							OUTRDA => SDATA,
							OUTFLAGA => OUTFLAGINST0
						);

	AL02: ORA00 PORT MAP(CLKO => CLK00,
							INFLAGO => OUTFLAGAC0,
							FUNCTO => FUNCT0,
							INRSO =>  INREGRS0,
							INRTO  => INREGRT0, 
							OUTRDO => SDATA,
							OUTFLAGO => OUTFLAGINST0
							);
	
	AL03: AC00 PORT MAP(CLKAC => CLK00,
							ENABLEAC => ENABLE0,
							INFLAGAC => OUTFLAGINST0,
							INAC => SDATA,
							OUTAC => OUTALU0,
							OUTFLAGAC => OUTFLAGAC0
						);

END A_TOPALU00;
