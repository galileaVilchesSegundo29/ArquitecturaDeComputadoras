LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY LCDCONTCONFIG00 IS
  PORT(
       CLKCC: IN STD_LOGIC;
       RESETCC: IN STD_LOGIC;
       INFLAGCC: IN STD_LOGIC;
       OUTCONTCC: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
       OUTFLAGCC: OUT STD_LOGIC);
END LCDCONTCONFIG00;

ARCHITECTURE A_LCDCONTCONFIG00 OF LCDCONTCONFIG00 IS
BEGIN
  PCONT: PROCESS(CLKCC)
  BEGIN
    IF (CLKCC'EVENT AND CLKCC = '1') THEN
      CASE RESETCC IS
        WHEN '0' =>
          OUTCONTCC <= (OTHERS => '0');
          OUTFLAGCC <= '0';
        WHEN '1' =>
          CASE INFLAGCC IS
            WHEN '0' =>
              OUTCONTCC <= OUTCONTCC + '1';
              OUTFLAGCC <= '1';
            WHEN '1' =>
              OUTCONTCC <= OUTCONTCC;
              OUTFLAGCC <= '0'; 
            WHEN OTHERS => NULL;
          END CASE;
        WHEN OTHERS => NULL;
      END CASE;
    END IF;
  END PROCESS PCONT;
END A_LCDCONTCONFIG00;

