LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY LCDMUX00 IS
  PORT(
       RESETM: IN STD_LOGIC;
       INFLAGCM: IN STD_LOGIC;
       INCOMMANDM: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
       INWORDM: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
       INRWCM: IN STD_LOGIC;
       INRSCM: IN STD_LOGIC;
       INENCM: IN STD_LOGIC;
       INRWDM: IN STD_LOGIC;
       INRSDM: IN STD_LOGIC;
       INENDM: IN STD_LOGIC;
       OUTWORDM: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
       OUTRWM: OUT STD_LOGIC;
       OUTRSM: OUT STD_LOGIC;
       OUTENM: OUT STD_LOGIC);
END LCDMUX00;

ARCHITECTURE A_LCDMUX00 OF LCDMUX00 IS
SIGNAL SCONTROL: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
SCONTROL <= (RESETM)&(INFLAGCM);
  WITH SCONTROL SELECT
     OUTWORDM <= INCOMMANDM WHEN "10",
                 INWORDM WHEN "11",
                 "00000000" WHEN OTHERS;

  WITH SCONTROL SELECT
     OUTRWM <= INRWCM WHEN "10",
               INRWDM WHEN "11",
               '0' WHEN OTHERS;

  WITH SCONTROL SELECT
     OUTRSM <= INRSCM WHEN "10",
               INRSDM WHEN "11",
               '0' WHEN OTHERS;

  WITH SCONTROL SELECT
     OUTENM <= INENCM WHEN "10",
               INENDM WHEN "11",
               '0' WHEN OTHERS;

END A_LCDMUX00;

