LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PACKAGELCD00 IS

  COMPONENT TOPDIV00
    PORT(
       CDIV0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
       CLK0: INOUT STD_LOGIC);
  END COMPONENT;
  
  COMPONENT LCDCONTCONFIG00
    PORT(
       CLKCC: IN STD_LOGIC;
       RESETCC: IN STD_LOGIC;
       INFLAGCC: IN STD_LOGIC;
       OUTCONTCC: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
       OUTFLAGCC: OUT STD_LOGIC);
  END COMPONENT;
  
  COMPONENT LCDCONFIG00
    PORT(
       CLKC: IN STD_LOGIC;
       RESETC: IN STD_LOGIC;
       INFLAGC: IN STD_LOGIC;
       INCONTC: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
       RWC: OUT STD_LOGIC;
       RSC: OUT STD_LOGIC;
       ENC: OUT STD_LOGIC;
       OUTCOMMANDC: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
       OUTFLAGC: OUT STD_LOGIC);
  END COMPONENT;
  
  COMPONENT LCDCONTDATA00
    PORT(
       CLKCD: IN STD_LOGIC;
       RESETCD: IN STD_LOGIC;
       INFLAGCD: IN STD_LOGIC;
       RWCD: OUT STD_LOGIC;
       RSCD: OUT STD_LOGIC;
       ENCD: OUT STD_LOGIC;
       OUTCONTCD: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0));
  END COMPONENT;
  
  COMPONENT LCDDATA00
  PORT(
       CLKD: IN STD_LOGIC;
       RESETD: IN STD_LOGIC;
       INFLAGD: IN STD_LOGIC;
       INCONTD: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
       OUTWORDD: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
  END COMPONENT;
  
  COMPONENT LCDMUX00
    PORT(
       RESETM: IN STD_LOGIC;
       INFLAGCM: IN STD_LOGIC;
       INCOMMANDM: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
       INRWCM: IN STD_LOGIC;
       INRSCM: IN STD_LOGIC;
       INENCM: IN STD_LOGIC;
       INWORDM: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
       INRWDM: IN STD_LOGIC;
       INRSDM: IN STD_LOGIC;
       INENDM: IN STD_LOGIC;
       OUTWORDM: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
       OUTRWM: OUT STD_LOGIC;
       OUTRSM: OUT STD_LOGIC;
       OUTENM: OUT STD_LOGIC);
  END COMPONENT;

END PACKAGELCD00;

