LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 
ENTITY EXSIGNO00 IS
   PORT(
        VECTOR_ENTRADA: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        VECTOR_SALIDA:  OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END EXSIGNO00 ;

ARCHITECTURE A_EXSIGNO00 OF EXSIGNO00  IS
SIGNAL VECTOR_AUXILIAR: STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN

    VECTOR_AUXILIAR <= "0000000000000000" & VECTOR_ENTRADA WHEN VECTOR_ENTRADA(15) = '0' 
    ELSE 
        "1111111111111111" & VECTOR_ENTRADA;
    VECTOR_SALIDA <= VECTOR_AUXILIAR; 

END A_EXSIGNO00;  

