LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY MUXSTACKB00 IS 
    PORT(
        RESETM, RWM: IN STD_LOGIC;
        INWORDCM, INWORDRM: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        OUTWORDM: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END MUXSTACKB00;

ARCHITECTURE A_MUXSTACKB00 OF MUXSTACKB00 IS
SIGNAL SCONTROLM: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
    SCONTROLM <= (RESETM)&(RWM);
    WITH SCONTROLM SELECT
        OUTWORDM <= INWORDCM WHEN "10",
                    INWORDRM WHEN "11",
                    "0000000" WHEN OTHERS;
END A_MUXSTACKB00;