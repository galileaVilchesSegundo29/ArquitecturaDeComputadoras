LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PACKAGEDIV00 IS

  COMPONENT OSC00
    PORT(OSC_INT: OUT STD_LOGIC);
  END COMPONENT;
  
  COMPONENT DIV00
    PORT(
       CLKDIV: IN STD_LOGIC;
     INDIV: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
       OUTDIV: INOUT STD_LOGIC);
  END COMPONENT;

END PACKAGEDIV00;

