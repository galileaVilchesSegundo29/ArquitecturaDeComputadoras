LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY MUXRAM00 IS 
    PORT(
        RESETM, RWM: IN STD_LOGIC;
        INWORDCM, INWORDRM: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        OUTWORDM: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END MUXRAM00;

ARCHITECTURE A_MUXRAM00 OF MUXRAM00 IS
SIGNAL SCONTROLM: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
    SCONTROLM <= (RESETM)&(RWM);
    WITH SCONTROLM SELECT
        OUTWORDM <= INWORDCM WHEN "10",
                    INWORDRM WHEN "11",
                    "0000000" WHEN OTHERS;
END A_MUXRAM00;