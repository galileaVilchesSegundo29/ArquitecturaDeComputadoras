LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGEBARRELRL00.ALL;

ENTITY TOPBARRELRL00 IS 
    PORT(
        CLK0: INOUT STD_LOGIC;
        CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        RESET0: IN STD_LOGIC;
        INS0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        INCON0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        OUTS0: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END TOPBARRELRL00;

ARCHITECTURE A_TOPBARRELRL00 OF TOPBARRELRL00 IS 
BEGIN
    SR00: topdiv00 PORT MAP(
        OSCOUT0 => CLK0,
        CDIV0 => CDIV00);
    SR01: barrelRL00 PORT MAP(
        CLKBRL => CLK0,
        INBRL => INS0,
        RESETBRL => RESET0,
        CONTROLBRL => INCON0,
        OUTBRL => OUTS0);
END A_TOPBARRELRL00;