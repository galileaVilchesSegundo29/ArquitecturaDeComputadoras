LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGEHA00 IS
    COMPONENT and00
        PORT(
            Aa, Ba: IN STD_LOGIC;
            Ya: OUT STD_LOGIC);
    END COMPONENT;

    COMPONENT xor00
        PORT(
            Ax, Bx: IN STD_LOGIC;
            Yx: OUT STD_LOGIC);
    END COMPONENT;
END PACKAGEHA00;
