LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGESHIFT00ALL IS
    COMPONENT topdiv00
        PORT(
            cdiv0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            oscout0: INOUT STD_LOGIC);
    END COMPONENT;

    COMPONENT shift00All
        PORT(
            CLKSFT, RESETSFT: IN STD_LOGIC;
            INRSSFT: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            INSELECTOR: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
            OUTRSSFT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
END PACKAGESHIFT00ALL;