LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGEDIV00 IS
    COMPONENT osc00
        PORT(
            OSC_INT: OUT STD_LOGIC);
    END COMPONENT;

    COMPONENT div00
        PORT(
            CLKDIV : IN STD_LOGIC;
            CDIV: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            OSCOUT: INOUT STD_LOGIC);
    END COMPONENT;
END PACKAGEDIV00;