LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY OSC00 IS
  PORT(OSC_INT: OUT STD_LOGIC);
END OSC00;

ARCHITECTURE A_OSC00 OF OSC00 IS
COMPONENT OSCH
   GENERIC (NOM_FREQ: STRING := "2.08");
   PORT ( STDBY :IN STD_LOGIC;
          OSC :OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE NOM_FREQ : STRING;
ATTRIBUTE NOM_FREQ OF OSCINST0 : LABEL IS "2.08";
BEGIN
   OSCINST0: OSCH
      GENERIC MAP ( NOM_FREQ => "2.08" )
      PORT MAP ( STDBY=> '0',
                OSC=> OSC_INT);
END A_OSC00;

