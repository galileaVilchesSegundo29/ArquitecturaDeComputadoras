LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY ORA00 IS
	PORT(
			CLKO: IN STD_LOGIC;
			INFLAGO: IN STD_LOGIC;
			FUNCTO: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			INRSO:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			INRTO:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);			
			OUTRDO:  OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			OUTFLAGO: OUT STD_LOGIC
		);
END ORA00;

ARCHITECTURE A_ORA00 OF ORA00 IS
BEGIN 
	POR: PROCESS(CLKO)
	VARIABLE AUX: BIT:='0';
	BEGIN 
		IF(CLKO'EVENT AND CLKO = '1') THEN
			IF (FUNCTO ="000001") THEN
				CASE INFLAGO IS
					WHEN '0'  =>
						OUTRDO <=(OTHERS => '0');
						OUTFLAGO <= '0';
					WHEN '1' =>
						IF (AUX ='0') THEN
							AUX:='1';
							OUTRDO <= INRSO OR INRTO;
							OUTFLAGO <='1';
						END IF;
					WHEN OTHERS => NULL;
				END CASE;
			ELSE
				AUX:='0';
				OUTRDO<=(OTHERS=>'Z');
				OUTFLAGO<='Z';
			END IF;
		END IF;
	END PROCESS POR;
END A_ORA00;
