LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGESHIFTRLR00 IS
    COMPONENT topdiv00
        PORT(
            cdiv0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            oscout0: INOUT STD_LOGIC);
    END COMPONENT;

    COMPONENT shiftrLR00
        PORT(
            CLKLR, RESETLR: IN STD_LOGIC;
            INRSLR: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            OUTRSLR: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
END PACKAGESHIFTRLR00;