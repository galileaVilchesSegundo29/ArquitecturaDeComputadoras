LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGEFA00 IS
    COMPONENT ha00
        PORT(
            A0, B0: IN STD_LOGIC;
            S0, C0: OUT STD_LOGIC);
    END COMPONENT;

    COMPONENT or00
        PORT(
            Ao, Bo: IN STD_LOGIC;
            Yo: OUT STD_LOGIC);
    END COMPONENT;
END PACKAGEFA00;