LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGEFA00.ALL;

ENTITY FA00 IS
    PORT(
        C00, A00, B00: IN STD_LOGIC;
        S00, C01: OUT STD_LOGIC);
END FA00;

ARCHITECTURE A_FA00 OF FA00 IS
SIGNAL SINT1:STD_LOGIC;
SIGNAL CINT1:STD_LOGIC;
SIGNAL CINT2:STD_LOGIC;
BEGIN 
    FA0: ha00 PORT MAP(
        A0 => A00,
        B0 => B00,
        S0 => SINT1,
        C0 => CINT1);
    FA01: ha00 PORT MAP(
        A0 => C00,
        B0 => SINT1,
        S0 => S00,
        C0 => CINT2);
    FA02: or00 PORT MAP(
        Ao => CINT2,
        Bo => CINT1,
        Yo => C01);
END A_FA00;