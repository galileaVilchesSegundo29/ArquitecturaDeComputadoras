LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;
USE PACKAGEROM00.ALL;

ENTITY TOPROM00 IS
    PORT(
        CLK0: INOUT STD_LOGIC;
        CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        RESET0: IN STD_LOGIC;
        CONT0: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        WORD0: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0);
        OUTTRANSIST0: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END TOPROM00;

ARCHITECTURE A_TOPROM00 OF TOPROM00 IS
BEGIN
    OUTTRANSIST0 <= "0001";

    RO00: topdiv00 PORT MAP(
            OSCOUT0 => CLK0,
            CDIV0 => CDIV00);
    
    RO02: contRead00 PORT MAP(
            CLKCR => CLK0,
            RESETCR => RESET0,
            OUTCONTCR => CONT0);

    RO03: rom00 PORT MAP(
            CLKRO => CLK0,
            RESETRO => RESET0,
            INDIRRO => CONT0,
            OUTWORDRO =>WORD0);
END A_TOPROM00;