LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PACKAGEWORD00 IS
    COMPONENT topdiv00
        PORT(
            cdiv0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            oscout0: INOUT STD_LOGIC);
    END COMPONENT;

    COMPONENT contring00 
        PORT(
            CLKS: IN STD_LOGIC;
            RESETS: IN STD_LOGIC;
            OUTS: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
    END COMPONENT;

    COMPONENT coder00
        PORT(
            INCONTC: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            OUTCODERC: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
    END COMPONENT;
END PACKAGEWORD00;