LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY LCDCONTDATA00 IS
  PORT(
       CLKCD: IN STD_LOGIC;
       RESETCD: IN STD_LOGIC;
       INFLAGCD: IN STD_LOGIC;
       RWCD: OUT STD_LOGIC;
       RSCD: OUT STD_LOGIC;
       ENCD: OUT STD_LOGIC;
       OUTCONTCD: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END LCDCONTDATA00;

ARCHITECTURE A_LCDCONTDATA00 OF LCDCONTDATA00 IS
SIGNAL SCONTROL: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
SCONTROL <= (RESETCD)&(INFLAGCD);
  PCD: PROCESS(CLKCD)
  VARIABLE AUX: BIT:='0';
  BEGIN
    IF (CLKCD'EVENT AND CLKCD = '1') THEN
      CASE SCONTROL IS
        WHEN "00" =>
          OUTCONTCD <= (OTHERS => '0');
        WHEN "11" =>
          IF ((OUTCONTCD < "01110")AND(AUX = '0')) THEN
              AUX:='1';
              OUTCONTCD <= OUTCONTCD + '1';
              RWCD <= '0';
              RSCD <= '1';
              ENCD <= '0';
          ELSIF ((OUTCONTCD < "01110")AND(AUX = '1')) THEN
              AUX:='0';
              OUTCONTCD <= OUTCONTCD;
              RWCD <= '0';
              RSCD <= '1';
              ENCD <= '1';
          END IF;
        WHEN OTHERS => NULL;
      END CASE;
    END IF;
  END PROCESS PCD;
END A_LCDCONTDATA00;

