LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGEBARREL00ALL.ALL;

ENTITY TOPBARREL00ALL IS 
    PORT(
        CLK0: INOUT STD_LOGIC;
        CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        RESET0: IN STD_LOGIC;
        INS0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        INSEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        INCON0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        OUTS0: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END TOPBARREL00ALL;

ARCHITECTURE A_TOPBARREL00ALL OF TOPBARREL00ALL IS 
BEGIN
    SR00: topdiv00 PORT MAP(
        OSCOUT0 => CLK0,
        CDIV0 => CDIV00);
    SR01: barrel00All PORT MAP(
        CLKBRL => CLK0,
        INBRL => INS0,
        INSELECTOR => INSEL,
        RESETBRL => RESET0,
        CONTROLBRL => INCON0,
        OUTBRL => OUTS0);
END A_TOPBARREL00ALL;