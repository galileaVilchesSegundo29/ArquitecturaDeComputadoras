LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGESHIFT00ALL.ALL;

ENTITY TOPSHIFT00ALL IS 
    PORT(
        CLK0: INOUT STD_LOGIC;
        CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        RESET0: IN STD_LOGIC;
        INS0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        INSEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        OUTS0: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END TOPSHIFT00ALL;

ARCHITECTURE A_TOPSHIFT00ALL OF TOPSHIFT00ALL IS 
BEGIN
    SR00: topdiv00 PORT MAP(
        OSCOUT0 => CLK0,
        CDIV0 => CDIV00);
    SR01: shift00All PORT MAP(
        CLKSFT => CLK0,
        INRSSFT => INS0,
        RESETSFT => RESET0,
        INSELECTOR => INSEL,
        OUTRSSFT => OUTS0);
END A_TOPSHIFT00ALL;