LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGESHIFTRLR00.ALL;

ENTITY TOPSHIFTRLR00 IS 
    PORT(
        CLK0: INOUT STD_LOGIC;
        CDIV00: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        RESET0: IN STD_LOGIC;
        INS0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        OUTS0: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END TOPSHIFTRLR00;

ARCHITECTURE A_TOPSHIFTRLR00 OF TOPSHIFTRLR00 IS 
BEGIN
    SR00: topdiv00 PORT MAP(
        OSCOUT0 => CLK0,
        CDIV0 => CDIV00);
    SR01: shiftrLR00 PORT MAP(
        CLKLR => CLK0,
        RESETLR => RESET0,
        INRSLR => INS0,
        OUTRSLR => OUTS0);
END A_TOPSHIFTRLR00;