LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE PACKAGEDIV00.ALL;

ENTITY TOPOSC00 IS
    PORT(
        OSCOUT0: INOUT STD_LOGIC;
        CDIV0: IN STD_LOGIC_VECTOR(4 DOWNTO 0)
    );
END TOPOSC00;

ARCHITECTURE A_TOPOSC00 OF TOPOSC00 IS
SIGNAL SCLK: STD_LOGIC;
BEGIN
    D00: OSC00 PORT MAP(
        OSC_INT => SCLK);

    D01: DIV00 PORT MAP(
        CLKDIV => SCLK,
        CDIV => CDIV0,
        OSCOUT => OSCOUT0);
END A_TOPOSC00;