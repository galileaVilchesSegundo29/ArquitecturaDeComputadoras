LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY MUXSTACKA00 IS 
    PORT(
        RESETM, RWM: IN STD_LOGIC;
        INWORDCM, INWORDRM: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        OUTWORDM: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END MUXSTACKA00;

ARCHITECTURE A_MUXSTACKA00 OF MUXSTACKA00 IS
SIGNAL SCONTROLM: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
    SCONTROLM <= (RESETM)&(RWM);
    WITH SCONTROLM SELECT
        OUTWORDM <= INWORDCM WHEN "10",
                    INWORDRM WHEN "11",
                    "0000000" WHEN OTHERS;
END A_MUXSTACKA00;