LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

PACKAGE PACKAGESHIFTRRL00 IS
    COMPONENT topdiv00
        PORT(
            cdiv0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            oscout0: INOUT STD_LOGIC);
    END COMPONENT;

    COMPONENT shiftrRL00
        PORT(
            CLKRL, RESETRL: IN STD_LOGIC;
            INRSRL: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            OUTRSRL: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
END PACKAGESHIFTRRL00;