LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY STACKA00 IS 
    PORT(
        CLKMRA: IN STD_LOGIC;
        RESETMRA: IN STD_LOGIC;
        RWMRA: IN STD_LOGIC;
        INDIRWMRA: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        INDIRRMRA: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        INWORDMRA: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        INFLAGMRA: IN STD_LOGIC;
        OUTWORDMRA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END STACKA00;

ARCHITECTURE A_STACKA00 OF STACKA00 IS
TYPE ARRAYSTACK IS ARRAY(0 TO 63) OF STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL WORDRAM: ARRAYSTACK;
SIGNAL SCONTROLM: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
    SCONTROLM <= (RESETMRA)&(RWMRA);
    PRAM: PROCESS(CLKMRA)
    BEGIN
        IF(CLKMRA'EVENT AND CLKMRA='1')THEN
            CASE SCONTROLM IS
                WHEN "10" =>
                    IF(INFLAGMRA = '1') THEN
                        WORDRAM(CONV_INTEGER(INDIRWMRA)) <= INWORDMRA;
                    END IF;
                WHEN "11" =>
                    OUTWORDMRA <= WORDRAM(CONV_INTEGER(INDIRRMRA));
                WHEN OTHERS => NULL;
            END CASE;
        END IF;
    END PROCESS PRAM;
END A_STACKA00;