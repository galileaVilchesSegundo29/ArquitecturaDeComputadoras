LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PACKAGEALU00 IS

	COMPONENT TOPDIV00
		PORT(
			CDIV0: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			CLK0: INOUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT ANDA00
		PORT(
			CLKA: IN STD_LOGIC;
			INFLAGA: IN STD_LOGIC;
			FUNCTA: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			INRSA:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			INRTA:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);			
			OUTRDA:  OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			OUTFLAGA: OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT ORA00
		PORT(
			CLKO: IN STD_LOGIC;
			INFLAGO: IN STD_LOGIC;
			FUNCTO: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			INRSO:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			INRTO:  IN STD_LOGIC_VECTOR (7 DOWNTO 0);			
			OUTRDO:  OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			OUTFLAGO: OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT AC00
		PORT(
			CLKAC: IN STD_LOGIC;
			ENABLEAC: IN STD_LOGIC;
			INFLAGAC: IN STD_LOGIC;
			INAC: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			OUTAC: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			OUTFLAGAC: OUT STD_LOGIC
		);
	END COMPONENT;
	
END PACKAGEALU00;
